module xor_gate(a,b,out);
output out;
input a,b;

      assign out = a^b;
endmodule