`include "mux4x1.v"

module mux4x1_str_tb();

    reg i0,i1,i2,i3,s1,s2;
    wire out;

  mux4x1_str DUT(out,i0,i1,i2,i3,s1,s2);

  initial 
  begin
   $monitor("At time %t,i0=(%0d),i1=(%0d),i2=(%0d),i3=(%0d),out=(%0d)",$time,i0,i1,i2,i3,out);
   $dumpfile("mux4x1_str_tb.vcd");
   $dumpvars(0, mux4x1_str_tb);

i0=0;i1=0;i2=0;i3=0;s1=0;s2=0;#1;
i0=0;i1=0;i2=0;i3=0;s1=0;s2=1;#1;
i0=0;i1=0;i2=0;i3=0;s1=1;s2=0;#1;
i0=0;i1=0;i2=0;i3=0;s1=1;s2=1;#1;

i0=0;i1=0;i2=0;i3=1;s1=0;s2=0;#1;
i0=0;i1=0;i2=0;i3=1;s1=0;s2=1;#1;
i0=0;i1=0;i2=0;i3=1;s1=1;s2=0;#1;
i0=0;i1=0;i2=0;i3=1;s1=1;s2=1;#1;

i0=0;i1=0;i2=1;i3=0;s1=0;s2=0;#1;
i0=0;i1=0;i2=1;i3=0;s1=0;s2=1;#1;
i0=0;i1=0;i2=1;i3=0;s1=1;s2=0;#1;
i0=0;i1=0;i2=1;i3=0;s1=1;s2=1;#1;

i0=0;i1=0;i2=1;i3=1;s1=0;s2=0;#1;
i0=0;i1=0;i2=1;i3=1;s1=0;s2=1;#1;
i0=0;i1=0;i2=1;i3=1;s1=1;s2=0;#1;
i0=0;i1=0;i2=1;i3=1;s1=1;s2=1;#1;

i0=0;i1=1;i2=0;i3=0;s1=0;s2=0;#1;
i0=0;i1=1;i2=0;i3=0;s1=0;s2=1;#1;
i0=0;i1=1;i2=0;i3=0;s1=1;s2=0;#1;
i0=0;i1=1;i2=0;i3=0;s1=1;s2=1;#1;

i0=0;i1=1;i2=0;i3=1;s1=0;s2=0;#1;
i0=0;i1=1;i2=0;i3=1;s1=0;s2=1;#1;
i0=0;i1=1;i2=0;i3=1;s1=1;s2=0;#1;
i0=0;i1=1;i2=0;i3=1;s1=1;s2=1;#1;

i0=0;i1=1;i2=1;i3=0;s1=0;s2=0;#1;
i0=0;i1=1;i2=1;i3=0;s1=0;s2=1;#1;
i0=0;i1=1;i2=1;i3=0;s1=1;s2=0;#1;
i0=0;i1=1;i2=1;i3=0;s1=1;s2=1;#1;

i0=0;i1=1;i2=1;i3=1;s1=0;s2=0;#1;
i0=0;i1=1;i2=1;i3=1;s1=0;s2=1;#1;
i0=0;i1=1;i2=1;i3=1;s1=1;s2=0;#1;
i0=0;i1=1;i2=1;i3=1;s1=1;s2=1;#1;

i0=1;i1=0;i2=0;i3=0;s1=0;s2=0;#1;
i0=1;i1=0;i2=0;i3=0;s1=0;s2=1;#1;
i0=1;i1=0;i2=0;i3=0;s1=1;s2=0;#1;
i0=1;i1=0;i2=0;i3=0;s1=1;s2=1;#1;

i0=1;i1=0;i2=0;i3=1;s1=0;s2=0;#1;
i0=1;i1=0;i2=0;i3=1;s1=0;s2=1;#1;
i0=1;i1=0;i2=0;i3=1;s1=1;s2=0;#1;
i0=1;i1=0;i2=0;i3=1;s1=1;s2=1;#1;

i0=1;i1=0;i2=1;i3=0;s1=0;s2=0;#1;
i0=1;i1=0;i2=1;i3=0;s1=0;s2=0;#1;
i0=1;i1=0;i2=1;i3=0;s1=0;s2=0;#1;
i0=1;i1=0;i2=1;i3=0;s1=0;s2=0;#1;

i0=1;i1=0;i2=1;i3=1;s1=0;s2=0;#1;
i0=1;i1=0;i2=1;i3=1;s1=0;s2=1;#1;
i0=1;i1=0;i2=1;i3=1;s1=1;s2=0;#1;
i0=1;i1=0;i2=1;i3=1;s1=1;s2=1;#1;

i0=1;i1=1;i2=0;i3=0;s1=0;s2=0;#1;
i0=1;i1=1;i2=0;i3=0;s1=0;s2=1;#1;
i0=1;i1=1;i2=0;i3=0;s1=1;s2=0;#1;
i0=1;i1=1;i2=0;i3=0;s1=1;s2=1;#1;

i0=1;i1=1;i2=0;i3=1;s1=0;s2=0;#1;
i0=1;i1=1;i2=0;i3=1;s1=0;s2=1;#1;
i0=1;i1=1;i2=0;i3=1;s1=1;s2=0;#1;
i0=1;i1=1;i2=0;i3=1;s1=1;s2=1;#1;

i0=1;i1=1;i2=1;i3=0;s1=0;s2=0;#1;
i0=1;i1=1;i2=1;i3=0;s1=0;s2=1;#1;
i0=1;i1=1;i2=1;i3=0;s1=1;s2=0;#1;
i0=1;i1=1;i2=1;i3=0;s1=1;s2=1;#1;

i0=1;i1=1;i2=1;i3=1;s1=0;s2=0;#1;
i0=1;i1=1;i2=1;i3=1;s1=0;s2=1;#1;
i0=1;i1=1;i2=1;i3=1;s1=1;s2=0;#1;
i0=1;i1=1;i2=1;i3=1;s1=1;s2=1;#1;

   end 
endmodule
   
     

