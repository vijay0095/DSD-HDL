module encoder_4x2(output y1,y0, input i3,i2,i1,i0);
or G1(y1,i3,i2);
or G2(y0,i3,i1);
endmodule
